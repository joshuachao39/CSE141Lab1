module InstROM #(parameter IW = 9, DW = 32)(
  input        [IW-1:0] InstAddress,	// address pointer
  output logic [DW-1:0] InstOut);

  logic [DW-1:0] inst_rom [2**IW];
  logic [8:0]    out      [2**IW];

  // load machine code program into instruction ROM
/*  initial begin
	$readmemb("C:/Users/riyang liu/Desktop/CSE-141L-lab4/CSE-141L-master/binary9.txt",out);
  end
*/
    for (genvar i = 0; i < out.size; i = i + 1) begin
        case (out[i])
            000000000 : inst_rom[i] = 0111_01_00000000000100000000000000;
            000000001 : inst_rom[i] = 0111_01_00010000001000000000000000;
            000000010 : inst_rom[i] = 0111_01_11100000001100000000000000;
            000000011 : inst_rom[i] = 0000_11_11010000000000000000000000;
            000000100 : inst_rom[i] = 0000_11_11000000000000000000000000;
            000000101 : inst_rom[i] = 0101_11_00000000000000110011000000;
            000000110 : inst_rom[i] = 0101_11_00010000000000110011000000;
            000000111 : inst_rom[i] = 0101_11_11100000000000110011000000;
            000001000 : inst_rom[i] = 0011_11_01000000000000000000000000;
            000001001 : inst_rom[i] = 0011_11_01110000000000000000000000;
            000001010 : inst_rom[i] = 0011_11_10010000000000000000000000;
            000001011 : inst_rom[i] = 0011_01_10010001000000010000000000;
            000001100 : inst_rom[i] = 0000_01_11111000000000000000000000;
            000001101 : inst_rom[i] = 0000_01_00100111000000000000000000;
            000001110 : inst_rom[i] = 0101_11_01000000100000100000000000;
            000001111 : inst_rom[i] = 0101_11_10010000000100010100000000;
            000010000 : inst_rom[i] = 1001_01_00010001000000010000000000;
            000010001 : inst_rom[i] = 0011_01_10010001000000010000000000;
            000010010 : inst_rom[i] = 0000_01_01000100000000010000000000;
            000010011 : inst_rom[i] = 0110_11_01000000100100001100000000;
            000010100 : inst_rom[i] = 0100_00_10100000010000000000000000;
            000010101 : inst_rom[i] = 0000_00_01110111101000000000000000;
            000010110 : inst_rom[i] = 0001_01_10001000000000000000000000;
            000010111 : inst_rom[i] = 0010_01_10110100111111110000000000;
            000011000 : inst_rom[i] = 0000_01_10111011000000010000000000;
            000011001 : inst_rom[i] = 0000_10_10100000100010110000000000;
            000011010 : inst_rom[i] = 1001_10_10111111111110100000000000;
            000011011 : inst_rom[i] = 0100_00_10111011101000000000000000;
            000011100 : inst_rom[i] = 0011_00_10110000101100000000000000;
            000011101 : inst_rom[i] = 1001_00_10111011101000000000000000;
            000011110 : inst_rom[i] = 0000_00_10001000101100000000000000;
            000011111 : inst_rom[i] = 0110_11_00110001000000010000000000;
            000100000 : inst_rom[i] = 0101_11_00110000100000110011000000;
            000100001 : inst_rom[i] = 0111_01_00010000001100000000000000;
            000100010 : inst_rom[i] = 0100_10_00000000000100110000000000;
            000100011 : inst_rom[i] = 0011_00_00000001000000000000000000;
            000100100 : inst_rom[i] = 1001_00_00000000001100000000000000;
            000100101 : inst_rom[i] = 0011_01_01000010100000000000000000;
            000100110 : inst_rom[i] = 1001_01_01000100000001110000000000;
            000100111 : inst_rom[i] = 0101_11_00000000000000101111000000;
            000101000 : inst_rom[i] = 0000_00_11001100001000000000000000;
            000101001 : inst_rom[i] = 0100_01_00100010000000010000000000;
            000101010 : inst_rom[i] = 0001_00_11011101111100000000000000;
            000101011 : inst_rom[i] = 0100_01_11111111000000010000000000;
            000101100 : inst_rom[i] = 0010_00_11111111010000000000000000;
            000101101 : inst_rom[i] = 0000_01_00110011000000010000000000;
            000101110 : inst_rom[i] = 0110_11_00110000100100100000000000;
            000101111 : inst_rom[i] = 0100_01_11111111000000010000000000;
            000110000 : inst_rom[i] = 0010_00_11111111010000000000000000;
            000110001 : inst_rom[i] = 0100_01_00100010000000010000000000;
            000110010 : inst_rom[i] = 0101_11_00000000000000101101000000;
            000110011 : inst_rom[i] = 1000_00_11010000010000000000000000;
            000110100 : inst_rom[i] = 1000_00_11000000010100000000000000;
            000110101 : inst_rom[i] = 1111_00_00000000000000000000000000;
            000110110 : inst_rom[i] = 0011_11_00000000000000000000000000;
            000110111 : inst_rom[i] = 0011_11_00010000000000000000000000;
            000111000 : inst_rom[i] = 0011_11_00100000000000000000000000;
            000111001 : inst_rom[i] = 0011_11_00110000000000000000000000;
            000111010 : inst_rom[i] = 0011_11_01000000000000000000000000;
            000111011 : inst_rom[i] = 0011_11_01010000000000000000000000;
            000111100 : inst_rom[i] = 0011_11_01100000000000000000000000;
            000111101 : inst_rom[i] = 0000_11_00000010000000000000000000;
            000111110 : inst_rom[i] = 0111_01_01000000010000000000000000;
            000111111 : inst_rom[i] = 0011_01_01000100000011110000000000;
            001000000 : inst_rom[i] = 0100_01_01000100000001000000000000;
            001000001 : inst_rom[i] = 0101_11_00000110000001010001000000;
            001000010 : inst_rom[i] = 0111_00_01010000000000000000000000;
            001000011 : inst_rom[i] = 0011_01_01100101111100000000000000;
            001000100 : inst_rom[i] = 0101_11_00010000010101001101000000;
            001000101 : inst_rom[i] = 0010_00_00110110010000000000000000;
            001000110 : inst_rom[i] = 0101_11_00110000000001001100000000;
            001000111 : inst_rom[i] = 0100_01_01010101000000010000000000;
            001001000 : inst_rom[i] = 0011_01_01100101111100000000000000;
            001001001 : inst_rom[i] = 0000_01_00010001000000010000000000;
            001001010 : inst_rom[i] = 0011_11_00110000000000000000000000;
            001001011 : inst_rom[i] = 0101_11_00110000000001000100000000;
            001001100 : inst_rom[i] = 0000_01_00100010000000010000000000;
            001001101 : inst_rom[i] = 0011_11_00010000000000000000000000;
            001001110 : inst_rom[i] = 0011_11_01100000000000000000000000;
            001001111 : inst_rom[i] = 0000_01_00000000000000010000000000;
            001010000 : inst_rom[i] = 0110_11_00000110000101000001000000;
            001010001 : inst_rom[i] = 1000_00_00100000011100000000000000;
            001010010 : inst_rom[i] = 1111_00_00000000000000000000000000;
            001010011 : inst_rom[i] = 0000_11_00010001010000000000000000;
            001010100 : inst_rom[i] = 0000_11_00100000000000000000000000;
            001010101 : inst_rom[i] = 0000_11_10000000000000000000000000;
            001010110 : inst_rom[i] = 0111_01_00111000000000000000000000;
            001010111 : inst_rom[i] = 0111_01_01001000100000000000000000;
            001011000 : inst_rom[i] = 0011_01_01010011010100000000000000;
            001011001 : inst_rom[i] = 0011_10_01000101000001100000000000;
            001011010 : inst_rom[i] = 0101_11_01010000000001011101000000;
            001011011 : inst_rom[i] = 0010_01_00110011111111110000000000;
            001011100 : inst_rom[i] = 0000_01_00110011000000010000000000;
            001011101 : inst_rom[i] = 0101_11_01100000000101100000000000;
            001011110 : inst_rom[i] = 0010_01_01000100111111110000000000;
            001011111 : inst_rom[i] = 0000_01_01000100000000010000000000;
            001100000 : inst_rom[i] = 0000_00_01110100001100000000000000;
            001100001 : inst_rom[i] = 0011_01_01110101010100000000000000;
            001100010 : inst_rom[i] = 0101_11_01010000000001100101000000;
            001100011 : inst_rom[i] = 0010_01_01110111111111110000000000;
            001100100 : inst_rom[i] = 0000_01_01110111000000010000000000;
            001100101 : inst_rom[i] = 0110_01_01111000011001110000000000;
            001100110 : inst_rom[i] = 0000_01_10000111000000000000000000;
            001100111 : inst_rom[i] = 0000_01_00100010000010000000000000;
            001101000 : inst_rom[i] = 0110_11_00101001000001010110000000;
            001101001 : inst_rom[i] = 0110_11_00010000000101110000000000;
            001101010 : inst_rom[i] = 0000_01_00010001111111110000000000;
            001101011 : inst_rom[i] = 0111_00_00110011000000000000000000;
            001101100 : inst_rom[i] = 0111_00_00110100000000000000000000;
            001101101 : inst_rom[i] = 0000_11_00100000000000000000000000;
            001101110 : inst_rom[i] = 0000_11_10100000000000000000000000;
            001101111 : inst_rom[i] = 0110_11_10100000000101011000000000;
            001110000 : inst_rom[i] = 1000_00_10000111111100000000000000;
            001110001 : inst_rom[i] = 1111_00_00000000000000000000000000;
            default   : inst_rom[i] = 1111_11_11111111111111111111111111;
        endcase
    end	  */
    // continuous combinational read output
    // change the pointer (from program counter) ==> change the output
    assign InstOut = inst_rom[InstAddress];
endmodule